xorGate