module not_(input a, output c);
				
assign c = !a;

				
endmodule